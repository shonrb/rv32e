module Execute (skid_buffer_port.upstream decoder);
endmodule
