parameter AHB_SLAVE_COUNT = 1;
parameter AHB_ADDR_MAP[AHB_SLAVE_COUNT-1] = '{
    default: 0
};

