export "DPI-C" task set_logging;

bit logging = 0;

task set_logging;
    logging = 1;
endtask



