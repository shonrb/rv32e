module Execute (input clock, input reset, skid_buffer_port.upstream decoder, bus_master.out bus);
    
endmodule
